-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus II License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 15.0.0 Build 145 04/22/2015 SJ Web Edition"
-- CREATED		"Tue Jan 23 18:01:52 2018"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY DE1_SOC_NIOS IS 
	PORT
	(
		CLOCK_50 :  IN  STD_LOGIC;
		DRAM_DQ :  INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		GPIO_00 :  IN  STD_LOGIC;
		GPIO_011 :  IN  STD_LOGIC;
		GPIO_128 :  IN  STD_LOGIC;
		GPIO_132 :  IN  STD_LOGIC;
		KEY :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		SW :  IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		DRAM_CLK :  OUT  STD_LOGIC;
		DRAM_CKE :  OUT  STD_LOGIC;
		DRAM_CS_N :  OUT  STD_LOGIC;
		DRAM_CAS_N :  OUT  STD_LOGIC;
		DRAM_RAS_N :  OUT  STD_LOGIC;
		DRAM_WE_N :  OUT  STD_LOGIC;
		DRAM_UDQM :  OUT  STD_LOGIC;
		DRAM_LDQM :  OUT  STD_LOGIC;
		VGA_HS :  OUT  STD_LOGIC;
		VGA_VS :  OUT  STD_LOGIC;
		VGA_BLANK_N :  OUT  STD_LOGIC;
		VGA_SYNC_N :  OUT  STD_LOGIC;
		VGA_CLK :  OUT  STD_LOGIC;
		DRAM_ADDR :  OUT  STD_LOGIC_VECTOR(12 DOWNTO 0);
		DRAM_BA :  OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		GPIO_05 :  OUT  STD_LOGIC;
		HEX0 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX1 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX2 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX3 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX4 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		HEX5 :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		LEDR :  OUT  STD_LOGIC_VECTOR(9 DOWNTO 0);
		VGA_B :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VGA_G :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		VGA_R :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END DE1_SOC_NIOS;

ARCHITECTURE bdf_type OF DE1_SOC_NIOS IS 

COMPONENT onchipm68xxio
	PORT(Clock_50Mhz : IN STD_LOGIC;
		 IOSelect_H : IN STD_LOGIC;
		 ByteSelect_L : IN STD_LOGIC;
		 WE_L : IN STD_LOGIC;
		 Reset_L : IN STD_LOGIC;
		 RS232_RxData : IN STD_LOGIC;
		 GPS_RxData : IN STD_LOGIC;
		 BlueTooth_RxData : IN STD_LOGIC;
		 TouchScreen_RxData : IN STD_LOGIC;
		 Address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 DataIn : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ACIA_IRQ : OUT STD_LOGIC;
		 RS232_TxData : OUT STD_LOGIC;
		 GPS_TxData : OUT STD_LOGIC;
		 BlueTooth_TxData : OUT STD_LOGIC;
		 TouchScreen_TxData : OUT STD_LOGIC;
		 DataOut : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT hexdisplays
	PORT(Hex0_1 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Hex2_3 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Hex4_5 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 HEX5 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT nios_ii_system
	PORT(CLOCK_50 : IN STD_LOGIC;
		 IO_acknowledge : IN STD_LOGIC;
		 IO_irq : IN STD_LOGIC;
		 DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 IO_read_data : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 KEY : IN STD_LOGIC_VECTOR(0 TO 0);
		 lcd_data : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Push_Buttons : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 DRAM_CLK : OUT STD_LOGIC;
		 DRAM_CKE : OUT STD_LOGIC;
		 DRAM_CS_N : OUT STD_LOGIC;
		 DRAM_CAS_N : OUT STD_LOGIC;
		 DRAM_RAS_N : OUT STD_LOGIC;
		 DRAM_WE_N : OUT STD_LOGIC;
		 DRAM_UDQM : OUT STD_LOGIC;
		 DRAM_LDQM : OUT STD_LOGIC;
		 IO_bus_enable : OUT STD_LOGIC;
		 IO_rw : OUT STD_LOGIC;
		 lcd_RS : OUT STD_LOGIC;
		 lcd_RW : OUT STD_LOGIC;
		 lcd_EN : OUT STD_LOGIC;
		 lcd_ON : OUT STD_LOGIC;
		 lcd_BLON : OUT STD_LOGIC;
		 DRAM_ADDR : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
		 DRAM_BA : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 Hex0_1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Hex2_3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 Hex4_5 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 IO_address : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 IO_byte_enable : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 IO_write_data : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT graphics_and_video_controller
	PORT(Reset_L : IN STD_LOGIC;
		 Clock_50Mhz : IN STD_LOGIC;
		 IOEnable_L : IN STD_LOGIC;
		 UpperByteSelect_L : IN STD_LOGIC;
		 LowerByteSelect_L : IN STD_LOGIC;
		 WriteEnable_L : IN STD_LOGIC;
		 GraphicsCS_L : IN STD_LOGIC;
		 Address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 DataIn : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 VGA_CLK : OUT STD_LOGIC;
		 VGA_HS : OUT STD_LOGIC;
		 VGA_VS : OUT STD_LOGIC;
		 VGA_BLANK_N : OUT STD_LOGIC;
		 DataOut : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 VGA_B : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VGA_G : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 VGA_R : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	gpio_10 :  STD_LOGIC;
SIGNAL	gpio_11 :  STD_LOGIC;
SIGNAL	gpio_111 :  STD_LOGIC;
SIGNAL	gpio_113 :  STD_LOGIC;
SIGNAL	gpio_115 :  STD_LOGIC;
SIGNAL	gpio_12 :  STD_LOGIC;
SIGNAL	GPIO_126 :  STD_LOGIC;
SIGNAL	gpio_13 :  STD_LOGIC;
SIGNAL	GPIO_134 :  STD_LOGIC;
SIGNAL	gpio_14 :  STD_LOGIC;
SIGNAL	gpio_15 :  STD_LOGIC;
SIGNAL	gpio_16 :  STD_LOGIC;
SIGNAL	gpio_17 :  STD_LOGIC;
SIGNAL	GPIO_ALTERA_SYNTHESIZED0 :  STD_LOGIC_VECTOR(11 DOWNTO 10);
SIGNAL	IO_byte_enable :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	IO_read_data :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	IO_write_data :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	DFF_inst14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;

SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN 
VGA_SYNC_N <= '0';
SYNTHESIZED_WIRE_7 <= '1';
SYNTHESIZED_WIRE_9 <= '1';

GDFX_TEMP_SIGNAL_0 <= (gpio_17 & gpio_16 & gpio_15 & gpio_14 & gpio_13 & gpio_12 & gpio_11 & gpio_10);


b2v_inst : onchipm68xxio
PORT MAP(Clock_50Mhz => CLOCK_50,
		 IOSelect_H => SYNTHESIZED_WIRE_18,
		 ByteSelect_L => SYNTHESIZED_WIRE_1,
		 WE_L => gpio_115,
		 Reset_L => SYNTHESIZED_WIRE_2,
		 RS232_RxData => GPIO_00,
		 GPS_RxData => GPIO_128,
		 BlueTooth_RxData => GPIO_132,
		 TouchScreen_RxData => GPIO_ALTERA_SYNTHESIZED0(11),
		 Address => SYNTHESIZED_WIRE_19,
		 DataIn => IO_write_data(7 DOWNTO 0),
		 ACIA_IRQ => SYNTHESIZED_WIRE_11,
		 RS232_TxData => GPIO_05,
		 TouchScreen_TxData => GPIO_ALTERA_SYNTHESIZED0(10),
		 DataOut => IO_read_data(7 DOWNTO 0));


b2v_inst1 : hexdisplays
PORT MAP(Hex0_1 => SYNTHESIZED_WIRE_4,
		 Hex2_3 => SYNTHESIZED_WIRE_5,
		 Hex4_5 => SYNTHESIZED_WIRE_6,
		 HEX0 => HEX0,
		 HEX1 => HEX1,
		 HEX2 => HEX2,
		 HEX3 => HEX3,
		 HEX4 => HEX4,
		 HEX5 => HEX5);


PROCESS(CLOCK_50,SYNTHESIZED_WIRE_7,SYNTHESIZED_WIRE_9)
BEGIN
IF (SYNTHESIZED_WIRE_7 = '0') THEN
	DFF_inst14 <= '0';
ELSIF (SYNTHESIZED_WIRE_9 = '0') THEN
	DFF_inst14 <= '1';
ELSIF (RISING_EDGE(CLOCK_50)) THEN
	DFF_inst14 <= SYNTHESIZED_WIRE_18;
END IF;
END PROCESS;





SYNTHESIZED_WIRE_20 <= NOT(SYNTHESIZED_WIRE_18);



SYNTHESIZED_WIRE_14 <= NOT(IO_byte_enable(0));



b2v_inst3 : nios_ii_system
PORT MAP(CLOCK_50 => CLOCK_50,
		 IO_acknowledge => DFF_inst14,
		 IO_irq => SYNTHESIZED_WIRE_11,
		 DRAM_DQ => DRAM_DQ,
		 IO_read_data => IO_read_data,
		 KEY(0) => KEY(0),
		 lcd_data => GDFX_TEMP_SIGNAL_0,
		 Push_Buttons => KEY(3 DOWNTO 1),
		 SW => SW,
		 DRAM_CLK => DRAM_CLK,
		 DRAM_CKE => DRAM_CKE,
		 DRAM_CS_N => DRAM_CS_N,
		 DRAM_CAS_N => DRAM_CAS_N,
		 DRAM_RAS_N => DRAM_RAS_N,
		 DRAM_WE_N => DRAM_WE_N,
		 DRAM_UDQM => DRAM_UDQM,
		 DRAM_LDQM => DRAM_LDQM,
		 IO_bus_enable => SYNTHESIZED_WIRE_18,
		 IO_rw => SYNTHESIZED_WIRE_15,
		 lcd_RW => gpio_115,
		 DRAM_ADDR => DRAM_ADDR,
		 DRAM_BA => DRAM_BA,
		 Hex0_1 => SYNTHESIZED_WIRE_4,
		 Hex2_3 => SYNTHESIZED_WIRE_5,
		 Hex4_5 => SYNTHESIZED_WIRE_6,
		 IO_address => SYNTHESIZED_WIRE_19,
		 IO_byte_enable => IO_byte_enable,
		 IO_write_data => IO_write_data,
		 LEDR => LEDR);


SYNTHESIZED_WIRE_13 <= NOT(IO_byte_enable(1));



SYNTHESIZED_WIRE_1 <= NOT(IO_byte_enable(0));



b2v_inst4 : graphics_and_video_controller
PORT MAP(Reset_L => KEY(0),
		 Clock_50Mhz => CLOCK_50,
		 IOEnable_L => SYNTHESIZED_WIRE_20,
		 UpperByteSelect_L => SYNTHESIZED_WIRE_13,
		 LowerByteSelect_L => SYNTHESIZED_WIRE_14,
		 WriteEnable_L => SYNTHESIZED_WIRE_15,
		 GraphicsCS_L => SYNTHESIZED_WIRE_20,
		 Address => SYNTHESIZED_WIRE_19,
		 DataIn => IO_write_data,
		 VGA_CLK => VGA_CLK,
		 VGA_HS => VGA_HS,
		 VGA_VS => VGA_VS,
		 VGA_BLANK_N => VGA_BLANK_N,
		 DataOut => IO_read_data,
		 VGA_B => VGA_B,
		 VGA_G => VGA_G,
		 VGA_R => VGA_R);


SYNTHESIZED_WIRE_2 <= NOT(KEY(0));



GPIO_ALTERA_SYNTHESIZED0(11) <= GPIO_011;
END bdf_type;